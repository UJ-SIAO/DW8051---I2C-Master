module HW3();


endmodule